module I2s{
    output  
}